// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Please do not spread this code without permission
module sram_128b_w2048 (CLK, D, Q, CEN, WEN, A);

  input  CLK;
  input  WEN;  // Write Enable (active low)
  input  CEN;  // Chip Enable (active low)
  input  [127:0] D;
  input  [10:0] A;
  output [127:0] Q;

  ////////// TECH INDEPENDENT ///////////
  // parameter num = 2048;

  // reg [127:0] memory [num-1:0];
  // reg [10:0] add_q = 0;
  // assign Q = memory[add_q];

  // integer i;
  // initial begin
  //   for (i = 0; i < num; i = i + 1) memory[i] = 128'b0;
  // end

  // always @ (posedge CLK) begin

  //  if (!CEN && WEN) // read 
  //     add_q <= A;
  //  if (!CEN && !WEN) // write
  //     memory[A] <= D; 

  // end

  ////////// TECH DEPENDENT -- IHP-SG13G2 ///////////
  // source: https://github.com/IHP-GmbH/IHP-Open-PDK/tree/main/ihp-sg13g2/libs.ref/sg13g2_sram
  genvar i;
  generate
    for (i = 0; i < 2; i = i+1) begin : gen_2048x64
      RM_IHPSG13_1P_2048x64_c2_bm_bist i_cut (
        .A_CLK (CLK),
        .A_DLY (1'b1),
        .A_ADDR(A),
        .A_BM  ({64{1'b1}}),
        .A_MEN (!CEN),
        .A_WEN (!WEN),
        .A_REN (WEN),
        .A_DIN (D[i*64 +: 64]),
        .A_DOUT(Q[i*64 +: 64]),
        .A_BIST_CLK (1'b0),
        .A_BIST_ADDR(11'd0),
        .A_BIST_DIN (64'd0),
        .A_BIST_BM  (64'd0),
        .A_BIST_MEN (1'b0),
        .A_BIST_WEN (1'b0),
        .A_BIST_REN (1'b0),
        .A_BIST_EN  (1'b0)
      );
    end
  endgenerate

endmodule
